

//My first project

module demo1(
  input a,
  output reg y
  
);
  
  assign y = a;
  
endmodule


