//My first project
//Author: Ryan Q. Nguyen

module demo1(
  input a,
  output reg y 
);
  
  assign y = a;
  
endmodule